// File: fifo_pkg.sv
package fifo_pkg;
  `include "uvm_macros.svh"
  import uvm_pkg::*;

  `include "fifo_seq_item.sv"
  `include "write_driver.sv"
  `include "read_driver.sv"
  `include "write_monitor.sv"
  `include "read_monitor.sv"
  `include "write_sequencer.sv"
  `include "read_sequencer.sv"
  `include "virtual_sequencer.sv"
  `include "write_sequence.sv"
  `include "read_seqwquence.sv"
  `include "virtual_sequence.sv"
  `include "write_agent.sv"
  `include "read_agent.sv"
  `include "fifo_coverage.sv"
  `include "fifo_scoreboard.sv"
  `include "fifo_env.sv"
  `include "base_test.sv"
endpackage
